`include "lib/defines.vh"

module cache_data(

);
endmodule