`include "lib/defines.vh"
module mem(
    input wire rst,

    input wire sel_rf_res,

    

);
endmodule 