`include "lib/defines.vh"

module cache_tag(

);
endmodule