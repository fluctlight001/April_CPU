`include "lib/defines.vh"
module dcache(
    input wire clk,
    input wire rst,

    input wire ex_pc
);



endmodule 