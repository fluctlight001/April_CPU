`include "defines.vh"
module decoder_6_64 (
    input wire [5:0] in,
    output reg [63:0] out
);
    always @ (*) begin
        case(in)
            6'd00:begin out=64'b0000000000000000000000000000000000000000000000000000000000000001; end
            6'd01:begin out=64'b0000000000000000000000000000000000000000000000000000000000000010; end
            6'd02:begin out=64'b0000000000000000000000000000000000000000000000000000000000000100; end
            6'd03:begin out=64'b0000000000000000000000000000000000000000000000000000000000001000; end
            6'd04:begin out=64'b0000000000000000000000000000000000000000000000000000000000010000; end
            6'd05:begin out=64'b0000000000000000000000000000000000000000000000000000000000100000; end
            6'd06:begin out=64'b0000000000000000000000000000000000000000000000000000000001000000; end
            6'd07:begin out=64'b0000000000000000000000000000000000000000000000000000000010000000; end
            6'd08:begin out=64'b0000000000000000000000000000000000000000000000000000000100000000; end
            6'd09:begin out=64'b0000000000000000000000000000000000000000000000000000001000000000; end
            6'd10:begin out=64'b0000000000000000000000000000000000000000000000000000010000000000; end
            6'd11:begin out=64'b0000000000000000000000000000000000000000000000000000100000000000; end
            6'd12:begin out=64'b0000000000000000000000000000000000000000000000000001000000000000; end
            6'd13:begin out=64'b0000000000000000000000000000000000000000000000000010000000000000; end
            6'd14:begin out=64'b0000000000000000000000000000000000000000000000000100000000000000; end
            6'd15:begin out=64'b0000000000000000000000000000000000000000000000001000000000000000; end
            6'd16:begin out=64'b0000000000000000000000000000000000000000000000010000000000000000; end
            6'd17:begin out=64'b0000000000000000000000000000000000000000000000100000000000000000; end
            6'd18:begin out=64'b0000000000000000000000000000000000000000000001000000000000000000; end
            6'd19:begin out=64'b0000000000000000000000000000000000000000000010000000000000000000; end
            6'd20:begin out=64'b0000000000000000000000000000000000000000000100000000000000000000; end
            6'd21:begin out=64'b0000000000000000000000000000000000000000001000000000000000000000; end
            6'd22:begin out=64'b0000000000000000000000000000000000000000010000000000000000000000; end
            6'd23:begin out=64'b0000000000000000000000000000000000000000100000000000000000000000; end
            6'd24:begin out=64'b0000000000000000000000000000000000000001000000000000000000000000; end
            6'd25:begin out=64'b0000000000000000000000000000000000000010000000000000000000000000; end
            6'd26:begin out=64'b0000000000000000000000000000000000000100000000000000000000000000; end
            6'd27:begin out=64'b0000000000000000000000000000000000001000000000000000000000000000; end
            6'd28:begin out=64'b0000000000000000000000000000000000010000000000000000000000000000; end
            6'd29:begin out=64'b0000000000000000000000000000000000100000000000000000000000000000; end
            6'd30:begin out=64'b0000000000000000000000000000000001000000000000000000000000000000; end
            6'd31:begin out=64'b0000000000000000000000000000000010000000000000000000000000000000; end
            6'd32:begin out=64'b0000000000000000000000000000000100000000000000000000000000000000; end
            6'd33:begin out=64'b0000000000000000000000000000001000000000000000000000000000000000; end
            6'd34:begin out=64'b0000000000000000000000000000010000000000000000000000000000000000; end
            6'd35:begin out=64'b0000000000000000000000000000100000000000000000000000000000000000; end
            6'd36:begin out=64'b0000000000000000000000000001000000000000000000000000000000000000; end
            6'd37:begin out=64'b0000000000000000000000000010000000000000000000000000000000000000; end
            6'd38:begin out=64'b0000000000000000000000000100000000000000000000000000000000000000; end
            6'd39:begin out=64'b0000000000000000000000001000000000000000000000000000000000000000; end
            6'd40:begin out=64'b0000000000000000000000010000000000000000000000000000000000000000; end
            6'd41:begin out=64'b0000000000000000000000100000000000000000000000000000000000000000; end
            6'd42:begin out=64'b0000000000000000000001000000000000000000000000000000000000000000; end
            6'd43:begin out=64'b0000000000000000000010000000000000000000000000000000000000000000; end
            6'd44:begin out=64'b0000000000000000000100000000000000000000000000000000000000000000; end
            6'd45:begin out=64'b0000000000000000001000000000000000000000000000000000000000000000; end
            6'd46:begin out=64'b0000000000000000010000000000000000000000000000000000000000000000; end
            6'd47:begin out=64'b0000000000000000100000000000000000000000000000000000000000000000; end
            6'd48:begin out=64'b0000000000000001000000000000000000000000000000000000000000000000; end
            6'd49:begin out=64'b0000000000000010000000000000000000000000000000000000000000000000; end
            6'd50:begin out=64'b0000000000000100000000000000000000000000000000000000000000000000; end
            6'd51:begin out=64'b0000000000001000000000000000000000000000000000000000000000000000; end
            6'd52:begin out=64'b0000000000010000000000000000000000000000000000000000000000000000; end
            6'd53:begin out=64'b0000000000100000000000000000000000000000000000000000000000000000; end
            6'd54:begin out=64'b0000000001000000000000000000000000000000000000000000000000000000; end
            6'd55:begin out=64'b0000000010000000000000000000000000000000000000000000000000000000; end
            6'd56:begin out=64'b0000000100000000000000000000000000000000000000000000000000000000; end
            6'd57:begin out=64'b0000001000000000000000000000000000000000000000000000000000000000; end
            6'd58:begin out=64'b0000010000000000000000000000000000000000000000000000000000000000; end
            6'd59:begin out=64'b0000100000000000000000000000000000000000000000000000000000000000; end
            6'd60:begin out=64'b0001000000000000000000000000000000000000000000000000000000000000; end
            6'd61:begin out=64'b0010000000000000000000000000000000000000000000000000000000000000; end
            6'd62:begin out=64'b0100000000000000000000000000000000000000000000000000000000000000; end
            6'd63:begin out=64'b1000000000000000000000000000000000000000000000000000000000000000; end   
            default:begin
                out=64'b0;
            end
        endcase
    end

endmodule 